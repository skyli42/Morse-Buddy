module MorseBuddy();

endmodule
